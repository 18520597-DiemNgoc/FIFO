library verilog;
use verilog.vl_types.all;
entity Compare_1bit is
    port(
        \Out\           : out    vl_logic;
        I0              : in     vl_logic;
        I1              : in     vl_logic
    );
end Compare_1bit;
